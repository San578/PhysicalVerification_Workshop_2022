**.subckt untitled in out
*.ipin in
*.opin out
x1 in GND out net1 inverter
V1 in GND PWL(0 0 20n 0 900n 1.8)
V2 net1 GND 1.8
**** begin user architecture code

.lib /usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt


.control
tran 1n 1u
plot V(in) V(out)
.endc

**** end user architecture code
**.ends

.include inverter.spice

.GLOBAL GND
** flattened .save nodes
.end
