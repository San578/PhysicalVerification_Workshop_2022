magic
tech sky130A
magscale 1 2
timestamp 1665753988
<< error_s >>
rect 508 2014 514 2020
rect 536 1986 542 2020
rect -50 1908 296 1978
rect -50 1644 -20 1908
rect 90 1880 324 1888
rect 162 1820 264 1846
rect 354 1820 456 1846
rect 190 1792 236 1818
rect 382 1792 428 1818
rect 286 1760 332 1770
rect 258 1732 360 1742
rect 190 1668 424 1672
rect -50 1572 396 1644
rect 536 1452 572 1748
rect 60 1076 288 1098
rect 88 1048 316 1070
rect 159 992 261 1002
rect 351 992 453 1002
rect 187 964 233 974
rect 379 964 425 974
rect 184 752 418 772
rect 156 724 390 744
<< pwell >>
rect -60 1908 296 1978
rect -60 1644 -20 1908
rect -60 1574 396 1644
rect -58 1572 396 1574
rect -66 1076 288 1146
rect -66 744 -22 1076
rect 536 986 572 1748
rect -66 680 390 744
rect -60 672 390 680
<< metal1 >>
rect 204 2268 404 2398
rect -26 2020 608 2268
rect -60 1908 296 1978
rect -60 1644 -20 1908
rect 536 1888 578 2020
rect 90 1820 578 1888
rect 536 1742 572 1748
rect 190 1668 572 1742
rect -60 1638 396 1644
rect -62 1572 396 1638
rect -718 1432 -518 1522
rect -62 1432 -26 1572
rect -718 1396 -26 1432
rect -718 1322 -518 1396
rect -62 1146 -26 1396
rect 536 1394 572 1668
rect 1056 1394 1256 1496
rect 536 1358 1256 1394
rect -66 1076 288 1146
rect -66 744 -22 1076
rect 536 1070 572 1358
rect 1056 1296 1256 1358
rect 88 992 576 1070
rect 536 986 572 992
rect 184 752 572 850
rect -66 680 390 744
rect -60 672 390 680
rect 458 622 568 752
rect -58 448 568 622
rect 138 328 338 448
use sky130_fd_pr__pfet_01v8_6LLYWG  XM2
timestamp 1665753988
transform 1 0 261 0 1 1771
box -311 -319 311 319
use sky130_fd_pr__nfet_01v8_RV7F6E  XM1
timestamp 1665753988
transform 1 0 258 0 1 907
box -311 -360 311 360
<< labels >>
flabel metal1 -718 1322 -518 1522 0 FreeSans 256 0 0 0 in
port 0 nsew
flabel metal1 1056 1296 1256 1496 0 FreeSans 256 0 0 0 out
port 3 nsew
flabel metal1 204 2198 404 2398 0 FreeSans 256 0 0 0 vdd
port 2 nsew
flabel metal1 138 328 338 528 0 FreeSans 256 0 0 0 vss
port 1 nsew
<< end >>
